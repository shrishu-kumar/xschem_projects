** sch_path: /home/shrishu/xschem_circuits/xor_sg_test.sch
**.subckt xor_sg_test
x1 vcc v1 vout v2 GND xor_sg
vcc vcc GND 1.8
V1 v1 GND pulse(0 1.8 0ns 0ns 0ns 5ns 10ns)
V2 v2 GND pulse(0 1.8 0ns 0ns 0ns 10ns 20ns)
**** begin user architecture code

.lib /home/shrishu/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 0.1n 80ns
.save all

**** end user architecture code
**.ends

* expanding   symbol:  xor_sg.sym # of pins=5
** sym_path: /home/shrishu/xschem_circuits/xor_sg.sym
** sch_path: /home/shrishu/xschem_circuits/xor_sg.sch
.subckt xor_sg vcc v1 vout v2 gnd
*.ipin vcc
*.opin vout
*.ipin v1
*.ipin v2
*.ipin gnd
x2 vcc v1 net2 net1 gnd Nand_Cmos
x3 vcc net2 vout net3 gnd Nand_Cmos
x4 vcc net1 net3 v2 gnd Nand_Cmos
x1 vcc v1 net1 v2 gnd Nand_Cmos
.ends


* expanding   symbol:  xschem_circuits/Nand_Cmos.sym # of pins=5
** sym_path: /home/shrishu/xschem_circuits/Nand_Cmos.sym
** sch_path: /home/shrishu/xschem_circuits/Nand_Cmos.sch
.subckt Nand_Cmos VDD A out B gnd
*.ipin B
*.ipin A
*.ipin VDD
*.ipin gnd
*.opin out
XM2 net2 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 A net1 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 B gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
C1 out gnd 0.12p m=1
R1 out net2 40 m=1
.ends

.GLOBAL GND
.end
