magic
tech sky130A
timestamp 1710978170
<< nwell >>
rect 55 15 200 195
<< nmos >>
rect 120 -65 135 -20
<< pmos >>
rect 120 35 135 95
<< ndiff >>
rect 75 -25 120 -20
rect 75 -60 85 -25
rect 105 -60 120 -25
rect 75 -65 120 -60
rect 135 -25 180 -20
rect 135 -60 150 -25
rect 170 -60 180 -25
rect 135 -65 180 -60
<< pdiff >>
rect 75 90 120 95
rect 75 40 85 90
rect 105 40 120 90
rect 75 35 120 40
rect 135 90 180 95
rect 135 40 150 90
rect 170 40 180 90
rect 135 35 180 40
<< ndiffc >>
rect 85 -60 105 -25
rect 150 -60 170 -25
<< pdiffc >>
rect 85 40 105 90
rect 150 40 170 90
<< psubdiff >>
rect 95 -110 160 -95
rect 95 -130 110 -110
rect 145 -130 160 -110
rect 95 -135 160 -130
<< nsubdiff >>
rect 80 160 165 170
rect 80 140 95 160
rect 145 140 165 160
rect 80 130 165 140
<< psubdiffcont >>
rect 110 -130 145 -110
<< nsubdiffcont >>
rect 95 140 145 160
<< poly >>
rect 120 95 135 115
rect 120 -20 135 35
rect 120 -85 135 -65
<< locali >>
rect 80 160 165 170
rect 80 140 95 160
rect 145 140 165 160
rect 80 130 165 140
rect 75 90 115 95
rect 75 40 85 90
rect 105 40 115 90
rect 75 35 115 40
rect 140 90 180 95
rect 140 40 150 90
rect 170 40 180 90
rect 140 35 180 40
rect 75 -25 115 -20
rect 75 -60 85 -25
rect 105 -60 115 -25
rect 75 -65 115 -60
rect 140 -25 180 -20
rect 140 -60 150 -25
rect 170 -60 180 -25
rect 140 -65 180 -60
rect 95 -110 160 -95
rect 95 -130 110 -110
rect 145 -130 160 -110
rect 95 -135 160 -130
<< end >>
