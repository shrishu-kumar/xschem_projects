** sch_path: /home/shrishu/xschem_circuits/INV_test.sch
**.subckt INV_test
x1 vcc v1 vout GND INVERTER
V1 v1 GND 0
V2 vcc GND 1.8
**** begin user architecture code

.lib /home/shrishu/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.dc v1 0 1.8 1m
.save all
.end

**** end user architecture code
**.ends

* expanding   symbol:  xschem_circuits/INVERTER.sym # of pins=4
** sym_path: /home/shrishu/xschem_circuits/INVERTER.sym
** sch_path: /home/shrishu/xschem_circuits/INVERTER.sch
.subckt INVERTER VDD VIN VOUT GND
*.ipin VIN
*.ipin VDD
*.ipin GND
*.opin VOUT
XM1 VOUT VIN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VOUT VIN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
